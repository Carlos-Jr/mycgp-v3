module top(pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16, po0, po1, po2, po3, po4, po5, po6, po7, po8);
  input pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8;
  wire n18, n19, n20, n21, n22, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34, n35, n36, n37, n38, n39, n40, n42, n43, n44, n45, n46, n47, n48, n49, n51, n52, n53, n54, n55, n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70, n71, n72, n73, n74, n75, n76, n78, n79, n80, n81, n82, n83, n84, n85, n87, n88;
  assign n18 = ~pi0 & pi8;
  assign n19 = pi0 & ~pi8;
  assign n20 = ~n18 & ~n19;
  assign n21 = pi16 & n20;
  assign n22 = ~pi16 & ~n20;
  assign po0 = n21 | n22;
  assign n24 = ~pi1 & pi9;
  assign n25 = pi1 & ~pi9;
  assign n26 = ~n24 & ~n25;
  assign n27 = pi16 & ~n20;
  assign n28 = pi0 & pi8;
  assign n29 = ~n27 & ~n28;
  assign n30 = n26 & ~n29;
  assign n31 = ~n26 & n29;
  assign po1 = n30 | n31;
  assign n33 = ~pi2 & pi10;
  assign n34 = pi2 & ~pi10;
  assign n35 = ~n33 & ~n34;
  assign n36 = ~n26 & ~n29;
  assign n37 = pi1 & pi9;
  assign n38 = ~n36 & ~n37;
  assign n39 = n35 & ~n38;
  assign n40 = ~n35 & n38;
  assign po2 = n39 | n40;
  assign n42 = ~pi3 & pi11;
  assign n43 = pi3 & ~pi11;
  assign n44 = ~n42 & ~n43;
  assign n45 = ~n35 & ~n38;
  assign n46 = pi2 & pi10;
  assign n47 = ~n45 & ~n46;
  assign n48 = n44 & ~n47;
  assign n49 = ~n44 & n47;
  assign po3 = n48 | n49;
  assign n51 = ~pi4 & pi12;
  assign n52 = pi4 & ~pi12;
  assign n53 = ~n51 & ~n52;
  assign n54 = ~n44 & ~n47;
  assign n55 = pi3 & pi11;
  assign n56 = ~n54 & ~n55;
  assign n57 = n53 & ~n56;
  assign n58 = ~n53 & n56;
  assign po4 = n57 | n58;
  assign n60 = ~pi5 & pi13;
  assign n61 = pi5 & ~pi13;
  assign n62 = ~n60 & ~n61;
  assign n63 = ~n53 & ~n56;
  assign n64 = pi4 & pi12;
  assign n65 = ~n63 & ~n64;
  assign n66 = n62 & ~n65;
  assign n67 = ~n62 & n65;
  assign po5 = n66 | n67;
  assign n69 = ~pi6 & pi14;
  assign n70 = pi6 & ~pi14;
  assign n71 = ~n69 & ~n70;
  assign n72 = ~n62 & ~n65;
  assign n73 = pi5 & pi13;
  assign n74 = ~n72 & ~n73;
  assign n75 = n71 & ~n74;
  assign n76 = ~n71 & n74;
  assign po6 = n75 | n76;
  assign n78 = ~pi7 & pi15;
  assign n79 = pi7 & ~pi15;
  assign n80 = ~n78 & ~n79;
  assign n81 = ~n71 & ~n74;
  assign n82 = pi6 & pi14;
  assign n83 = ~n81 & ~n82;
  assign n84 = n80 & ~n83;
  assign n85 = ~n80 & n83;
  assign po7 = n84 | n85;
  assign n87 = ~n80 & ~n83;
  assign n88 = pi7 & pi15;
  assign po8 = n87 | n88;
endmodule
